module mux_template(
  
)
  endmodule
